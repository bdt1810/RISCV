`timescale 1ns / 1ps
module tb_RISCV;
	reg clk;
	initial 
	begin
		clk=0;
		forever #200
		clk= ~clk;
	end
	RISCV RISCV(clk);

endmodule
